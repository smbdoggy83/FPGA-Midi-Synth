module MidiNoteNumberToSampleTicks_verilog(
	input [7:0] midiNoteNumber,
	output reg [23:0] noteSampleTicks
);

always @(midiNoteNumber)
begin
	case (midiNoteNumber)
		8'h00: noteSampleTicks <= 24'd23889;  // 0
		8'h01: noteSampleTicks <= 24'd22548;  // 1
		8'h02: noteSampleTicks <= 24'd21282;  // 2
		8'h03: noteSampleTicks <= 24'd20088;  // 3
		8'h04: noteSampleTicks <= 24'd18960;  // 4
		8'h05: noteSampleTicks <= 24'd17896;  // 5
		8'h06: noteSampleTicks <= 24'd16892;  // 6
		8'h07: noteSampleTicks <= 24'd15944;  // 7
		8'h08: noteSampleTicks <= 24'd15049;  // 8
		8'h09: noteSampleTicks <= 24'd14204;  // 9
		8'h0A: noteSampleTicks <= 24'd13407;  // 10
		8'h0B: noteSampleTicks <= 24'd12654;  // 11
		8'h0C: noteSampleTicks <= 24'd11944;  // 12
		8'h0D: noteSampleTicks <= 24'd11274;  // 13
		8'h0E: noteSampleTicks <= 24'd10641;  // 14
		8'h0F: noteSampleTicks <= 24'd10044;  // 15
		8'h10: noteSampleTicks <= 24'd9480;  // 16
		8'h11: noteSampleTicks <= 24'd8948;  // 17
		8'h12: noteSampleTicks <= 24'd8446;  // 18
		8'h13: noteSampleTicks <= 24'd7972;  // 19
		8'h14: noteSampleTicks <= 24'd7524;  // 20
		8'h15: noteSampleTicks <= 24'd7102;  // 21
		8'h16: noteSampleTicks <= 24'd6703;  // 22
		8'h17: noteSampleTicks <= 24'd6327;  // 23
		8'h18: noteSampleTicks <= 24'd5972;  // 24
		8'h19: noteSampleTicks <= 24'd5637;  // 25
		8'h1A: noteSampleTicks <= 24'd5320;  // 26
		8'h1B: noteSampleTicks <= 24'd5022;  // 27
		8'h1C: noteSampleTicks <= 24'd4740;  // 28
		8'h1D: noteSampleTicks <= 24'd4474;  // 29
		8'h1E: noteSampleTicks <= 24'd4223;  // 30
		8'h1F: noteSampleTicks <= 24'd3986;  // 31
		8'h20: noteSampleTicks <= 24'd3762;  // 32
		8'h21: noteSampleTicks <= 24'd3551;  // 33
		8'h22: noteSampleTicks <= 24'd3351;  // 34
		8'h23: noteSampleTicks <= 24'd3163;  // 35
		8'h24: noteSampleTicks <= 24'd2986;  // 36
		8'h25: noteSampleTicks <= 24'd2818;  // 37
		8'h26: noteSampleTicks <= 24'd2660;  // 38
		8'h27: noteSampleTicks <= 24'd2511;  // 39
		8'h28: noteSampleTicks <= 24'd2370;  // 40
		8'h29: noteSampleTicks <= 24'd2237;  // 41
		8'h2A: noteSampleTicks <= 24'd2111;  // 42
		8'h2B: noteSampleTicks <= 24'd1993;  // 43
		8'h2C: noteSampleTicks <= 24'd1881;  // 44
		8'h2D: noteSampleTicks <= 24'd1775;  // 45
		8'h2E: noteSampleTicks <= 24'd1675;  // 46
		8'h2F: noteSampleTicks <= 24'd1581;  // 47
		8'h30: noteSampleTicks <= 24'd1493;  // 48
		8'h31: noteSampleTicks <= 24'd1409;  // 49
		8'h32: noteSampleTicks <= 24'd1330;  // 50
		8'h33: noteSampleTicks <= 24'd1255;  // 51
		8'h34: noteSampleTicks <= 24'd1185;  // 52
		8'h35: noteSampleTicks <= 24'd1118;  // 53
		8'h36: noteSampleTicks <= 24'd1055;  // 54
		8'h37: noteSampleTicks <= 24'd996;  // 55
		8'h38: noteSampleTicks <= 24'd940;  // 56
		8'h39: noteSampleTicks <= 24'd887;  // 57
		8'h3A: noteSampleTicks <= 24'd837;  // 58
		8'h3B: noteSampleTicks <= 24'd790;  // 59
		8'h3C: noteSampleTicks <= 24'd746;  // 60
		8'h3D: noteSampleTicks <= 24'd704;  // 61
		8'h3E: noteSampleTicks <= 24'd665;  // 62
		8'h3F: noteSampleTicks <= 24'd627;  // 63
		8'h40: noteSampleTicks <= 24'd592;  // 64
		8'h41: noteSampleTicks <= 24'd559;  // 65
		8'h42: noteSampleTicks <= 24'd527;  // 66
		8'h43: noteSampleTicks <= 24'd498;  // 67
		8'h44: noteSampleTicks <= 24'd470;  // 68
		8'h45: noteSampleTicks <= 24'd443;  // 69
		8'h46: noteSampleTicks <= 24'd418;  // 70
		8'h47: noteSampleTicks <= 24'd395;  // 71
		8'h48: noteSampleTicks <= 24'd373;  // 72
		8'h49: noteSampleTicks <= 24'd352;  // 73
		8'h4A: noteSampleTicks <= 24'd332;  // 74
		8'h4B: noteSampleTicks <= 24'd313;  // 75
		8'h4C: noteSampleTicks <= 24'd296;  // 76
		8'h4D: noteSampleTicks <= 24'd279;  // 77
		8'h4E: noteSampleTicks <= 24'd263;  // 78
		8'h4F: noteSampleTicks <= 24'd249;  // 79
		8'h50: noteSampleTicks <= 24'd235;  // 80
		8'h51: noteSampleTicks <= 24'd221;  // 81
		8'h52: noteSampleTicks <= 24'd209;  // 82
		8'h53: noteSampleTicks <= 24'd197;  // 83
		8'h54: noteSampleTicks <= 24'd186;  // 84
		8'h55: noteSampleTicks <= 24'd176;  // 85
		8'h56: noteSampleTicks <= 24'd166;  // 86
		8'h57: noteSampleTicks <= 24'd156;  // 87
		8'h58: noteSampleTicks <= 24'd148;  // 88
		8'h59: noteSampleTicks <= 24'd139;  // 89
		8'h5A: noteSampleTicks <= 24'd131;  // 90
		8'h5B: noteSampleTicks <= 24'd124;  // 91
		8'h5C: noteSampleTicks <= 24'd117;  // 92
		8'h5D: noteSampleTicks <= 24'd110;  // 93
		8'h5E: noteSampleTicks <= 24'd104;  // 94
		8'h5F: noteSampleTicks <= 24'd98;  // 95
		8'h60: noteSampleTicks <= 24'd93;  // 96
		8'h61: noteSampleTicks <= 24'd88;  // 97
		8'h62: noteSampleTicks <= 24'd83;  // 98
		8'h63: noteSampleTicks <= 24'd78;  // 99
		8'h64: noteSampleTicks <= 24'd74;  // 100
		8'h65: noteSampleTicks <= 24'd69;  // 101
		8'h66: noteSampleTicks <= 24'd65;  // 102
		8'h67: noteSampleTicks <= 24'd62;  // 103
		8'h68: noteSampleTicks <= 24'd58;  // 104
		8'h69: noteSampleTicks <= 24'd55;  // 105
		8'h6A: noteSampleTicks <= 24'd52;  // 106
		8'h6B: noteSampleTicks <= 24'd49;  // 107
		8'h6C: noteSampleTicks <= 24'd46;  // 108
		8'h6D: noteSampleTicks <= 24'd44;  // 109
		8'h6E: noteSampleTicks <= 24'd41;  // 110
		8'h6F: noteSampleTicks <= 24'd39;  // 111
		8'h70: noteSampleTicks <= 24'd37;  // 112
		8'h71: noteSampleTicks <= 24'd34;  // 113
		8'h72: noteSampleTicks <= 24'd32;  // 114
		8'h73: noteSampleTicks <= 24'd31;  // 115
		8'h74: noteSampleTicks <= 24'd29;  // 116
		8'h75: noteSampleTicks <= 24'd27;  // 117
		8'h76: noteSampleTicks <= 24'd26;  // 118
		8'h77: noteSampleTicks <= 24'd24;  // 119
		8'h78: noteSampleTicks <= 24'd23;  // 120
		8'h79: noteSampleTicks <= 24'd22;  // 121
		8'h7A: noteSampleTicks <= 24'd20;  // 122
		8'h7B: noteSampleTicks <= 24'd19;  // 123
		8'h7C: noteSampleTicks <= 24'd18;  // 124
		8'h7D: noteSampleTicks <= 24'd17;  // 125
		8'h7E: noteSampleTicks <= 24'd16;  // 126
		8'h7F: noteSampleTicks <= 24'd15;  // 127

		default: noteSampleTicks <= 0;
	endcase
end

endmodule
