module Top_Level_ver(
	// Synth
	input CLOCK_50,
	input MIDI_RX, 
//	output reg I2S_BIT_CLOCK, // Not used
//	output reg I2S_SOUND_DATA, // Goes to i2sound instead of direct output
//	output reg I2S_LEFT_RIGHT_SELECT, // Not used
	output reg [9:0] LEDR,

	// i2sound
	input [3:0] KEY,
	output reg [6:0] HEX0,
	output reg [6:0] HEX1,
	input AUD_ADCDAT,				// Audio in (Physical)
	output reg AUD_DACDAT, 		// Audio Out
	output reg AUD_XCK,
	output reg FPGA_I2C_SCLK,
	inout FPGA_I2C_SDAT,

	// Other
	input [9:0] SW // Toggle Audio Source / Filter
);

wire isNoteOn;
wire [23:0] noteSampleTicks;
wire [7:0] modulationValue;

wire [9:0] ledr;
wire [6:0] hex0;
wire [6:0] hex1;
wire aud_dacdat;
wire aud_xck;

reg filter_in;
reg audio_in;

SoundModule soundmodule(CLOCK_50, MIDI_RX, i2s_bit_clock, i2s_sound_data, i2s_left_right_select, ledr); // Synthesizer itself
bandpass_leastPth_ver filter(CLOCK_50, 1'b1, 1'b0, filter_in, filter_out); // Bandpass Filter
DE10_Standard_i2sound i2sound(CLOCK_50, KEY, hex0, hex1, audio_in, aud_dacdat, aud_xck, fpga_i2c_sclk, FPGA_I2C_SDAT); // Audio In / Out


always @(posedge CLOCK_50)
begin
	LEDR <= ledr;
	HEX0 <= hex0;
	HEX1 <= hex1;
	AUD_DACDAT <= aud_dacdat; // audio output
	AUD_XCK <= aud_xck;
	FPGA_I2C_SCLK <= fpga_i2c_sclk;

	filter_in <= SW[0] ? i2s_sound_data : AUD_ADCDAT; // Switch 0 Controls if audio is from synth or from physical jack
	audio_in <= SW[1] ? filter_out : filter_in; // Switch 1 Controls if filter is enabled 	
end


endmodule


//=======================================================
//  This code is generated by Terasic System Builder
//=======================================================

module DE10_Standard_i2sound(

//	//////////// CLOCK //////////
//	input 		          		CLOCK2_50,
//	input 		          		CLOCK3_50,
//	input 		          		CLOCK4_50,
	input 		          		CLOCK_50,

	//////////// KEY //////////
	input 		     [3:0]		KEY,


//	output		     [9:0]		LEDR,

	//////////// Seg7 //////////
	output		     [6:0]		HEX0,
	output		     [6:0]		HEX1,
//	output		     [6:0]		HEX2,
//	output		     [6:0]		HEX3,
//	output		     [6:0]		HEX4,
//	output		     [6:0]		HEX5,

	//////////// Audio //////////
	input 		          		AUD_ADCDAT,
//	inout 		          		AUD_ADCLRCK,
//	inout 		          		AUD_BCLK,
	output		          		AUD_DACDAT,
//	inout 		          		AUD_DACLRCK,
	output		          		AUD_XCK,

	//////////// I2C for Audio and Video-In //////////
	output		          		FPGA_I2C_SCLK,
	inout 		          		FPGA_I2C_SDAT

);



///=======================================================
//  REG/WIRE declarations
//=======================================================
wire				CLK_1M;
wire			 	END;
wire			 	KEY0_EDGE;
wire	[23:0] 		AUD_I2C_DATA;
wire         		GO;
wire  	[3:0]  		level_vol;
wire [23:0] 	audio_out;
reg  [23:0]    audio_out_reg;

//=======================================================
//  Structural coding
//=======================================================
assign		LEDR = 10'h000;
assign		HEX1 = 7'h40;
assign		AUD_DACDAT = AUD_ADCDAT;

//KEY triggle - Takes in the button (key) and uses the clock to debounce it, returns a signal that just represents the pressing-in-edge of pressing the button
keytr			u3( 
	.clock(CLK_1M),
	.key0(KEY[0]),
	.rst_n(KEY[1]),
	
	.KEY0_EDGE(KEY0_EDGE)
	);

//I2C output data
CLOCK_500		u1(
	.CLOCK(CLOCK_50), //The Outputting Clock Signal is Connected to the CLOCK_50 Signal on the DE-10
	.rst_n(KEY[1]), // The Reset Signal is Connected to KEY1 on the DE-10					 
	.END(END), //Stopping the Process of Outputting the I2C Data to the I2S on the DE-10
	.KEY0_EDGE(KEY0_EDGE), //The Edge Signal for KEY0 is Connected to the Edge Signal for KEY0 on the DE-10
	
	.CLOCK_500(CLK_1M), //The Clock_500 Signal Outputting from the I2C is Connected to a 1MHz on the DE-10
	.GO(GO), //Process of Moving the I2C Serial Data             
	.CLOCK_2(AUD_XCK), //The Clock_2 Signal Outputting from the I2C is Connected to the Audio XCK Signal on the I2S in the DE-10
	.DATA(AUD_I2C_DATA), //The Data Signal Outputting from the I2C is Connected to the Audio I2C Data Signal on the I2S in the DE-10
	.level_vol(level_vol) //The Outputting Volume Level is Mapped to the I2C Volume Level on the DE-10
	);
					 
//i2c input controller
i2c				u2( 
	// Host Side
	.CLOCK(CLK_1M), //The Overall Clock Signal from the Controller is Connected to a 1MHz Clock on the DE-10
	.RESET(1'b1), //The Reset Signal from the Controller is Connected to the Value 1'b1 on the DE-10
	// I2C Side
	.I2C_SDAT(FPGA_I2C_SDAT), //The I2C Data Signal from the Controller is Connected to the FPGA I2C Data Signal for the Audio In of the I2S on the DE-10
	.I2C_DATA(AUD_I2C_DATA), //The 24 Bit I2C Serial Data from the Controller is Connected to the 24 Bit Audio I2C Data Signal for the I2S on the DE-10
	.I2C_SCLK(FPGA_I2C_SCLK), //The I2C Clock Signal from the Controller is Connected to the FPGA I2C Clock Signal for the Audio In of the I2S on the DE-10
	// Control Signals
	.GO(GO), //Process of Moving the I2C Serial Data
	.END(END) //Stopping the Process of Moving I2C Serial Data
	);
					 
HEX				u4(
	.hex(level_vol), 
	.hex_fps(HEX0) //Displays the Volume Level on the DE-10
	);

endmodule

module SoundModule(
	input CLOCK_50,
	input MIDI_RX,
	output reg I2S_BIT_CLOCK,
	output reg I2S_SOUND_DATA,
	output reg I2S_LEFT_RIGHT_SELECT,
	output reg [7:0] LEDR
);

wire i2sBitClock;
wire i2sSoundData;
wire i2sLeftRightSelect;

wire isNoteOn;
wire [23:0] noteSampleTicks;
wire [7:0] modulationValue;

MidiProcessor midiProcessor(CLOCK_50, MIDI_RX, isNoteOn, noteSampleTicks, modulationValue);
Synthesizer synthesizer(CLOCK_50, isNoteOn, noteSampleTicks, modulationValue, i2sBitClock, i2sSoundData, i2sLeftRightSelect);

always @(posedge CLOCK_50)
begin
	I2S_BIT_CLOCK <= i2sBitClock;
	I2S_SOUND_DATA <= i2sSoundData;
	I2S_LEFT_RIGHT_SELECT <= i2sLeftRightSelect;

	LEDR <= isNoteOn ? noteSampleTicks[7:0] : 8'h00;
end

endmodule

// -------------------------------------------------------------
//
// Module: bandpass_leastPth_ver
// Generated by MATLAB(R) 9.11 and Filter Design HDL Coder 3.1.10.
// Generated on: 2022-05-01 14:21:29
// -------------------------------------------------------------

// -------------------------------------------------------------
// HDL Code Generation Options:
//
// Name: bandpass_leastPth_ver
// TargetLanguage: Verilog
// TestBenchStimulus: step ramp chirp 
// GenerateHDLTestBench: off

// Filter Specifications:
//
// Sample Rate            : N/A (normalized frequency)
// Response               : Bandpass
// Specification          : Fst1,Fp1,Fp2,Fst2,Ast1,Ap,Ast2
// First Stopband Edge    : 0.35
// Second Stopband Atten. : 60 dB
// Passband Ripple        : 1 dB
// Second Passband Edge   : 0.55
// First Passband Edge    : 0.45
// Second Stopband Edge   : 0.65
// First Stopband Atten.  : 60 dB
// -------------------------------------------------------------

// -------------------------------------------------------------
// HDL Implementation    : Fully parallel
// Folding Factor        : 1
// -------------------------------------------------------------
// Filter Settings:
//
// Discrete-Time IIR Filter (real)
// -------------------------------
// Filter Structure    : Direct-Form II, Second-Order Sections
// Number of Sections  : 12
// Stable              : Yes
// Linear Phase        : No
// Arithmetic          : fixed
// Numerator           : s24,21 -> [-4 4)
// Denominator         : s24,22 -> [-2 2)
// Scale Values        : s24,34 -> [-4.882812e-04 4.882812e-04)
// Input               : s24,23 -> [-1 1)
// Section Input       : s24,28 -> [-3.125000e-02 3.125000e-02)
// Section Output      : s24,18 -> [-32 32)
// Output              : s24,18 -> [-32 32)
// State               : s24,23 -> [-1 1)
// Numerator Prod      : s48,44 -> [-8 8)
// Denominator Prod    : s48,45 -> [-4 4)
// Numerator Accum     : s40,34 -> [-32 32)
// Denominator Accum   : s40,35 -> [-16 16)
// Round Mode          : convergent
// Overflow Mode       : wrap
// Cast Before Sum     : true
// -------------------------------------------------------------




`timescale 1 ns / 1 ns

module bandpass_leastPth_ver
               (
                clk,
                clk_enable,
                reset,
                filter_in,
                filter_out
                );

  input   clk; 
  input   clk_enable; 
  input   reset; 
  input   signed [23:0] filter_in; //sfix24_En23
  output  signed [23:0] filter_out; //sfix24_En18

////////////////////////////////////////////////////////////////
//Module Architecture: bandpass_leastPth_ver
////////////////////////////////////////////////////////////////
  // Local Functions
  // Type Definitions
  // Constants
  parameter signed [23:0] scaleconst1 = 24'b101011011110111000111100; //sfix24_En34
  parameter signed [23:0] coeff_b1_section1 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section1 = 24'b110100011011000001111000; //sfix24_En21
  parameter signed [23:0] coeff_b3_section1 = 24'b000011100101000000000000; //sfix24_En21
  parameter signed [23:0] coeff_a2_section1 = 24'b100001111110000111100011; //sfix24_En22
  parameter signed [23:0] coeff_a3_section1 = 24'b001110011101001010101001; //sfix24_En22
  parameter signed [23:0] coeff_b1_section2 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section2 = 24'b000100100110001000011001; //sfix24_En21
  parameter signed [23:0] coeff_b3_section2 = 24'b000000001100011011110110; //sfix24_En21
  parameter signed [23:0] coeff_a2_section2 = 24'b100001011111010111011100; //sfix24_En22
  parameter signed [23:0] coeff_a3_section2 = 24'b001111101000010110000110; //sfix24_En22
  parameter signed [23:0] coeff_b1_section3 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section3 = 24'b110000110101001110110011; //sfix24_En21
  parameter signed [23:0] coeff_b3_section3 = 24'b000111111111100111000111; //sfix24_En21
  parameter signed [23:0] coeff_a2_section3 = 24'b100010000010100101100000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section3 = 24'b001110110011110111000000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section4 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section4 = 24'b110111010000001101100010; //sfix24_En21
  parameter signed [23:0] coeff_b3_section4 = 24'b000000110000001010010100; //sfix24_En21
  parameter signed [23:0] coeff_a2_section4 = 24'b100001000101000011101110; //sfix24_En22
  parameter signed [23:0] coeff_a3_section4 = 24'b001111000101010011101000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section5 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section5 = 24'b111110111101010001101111; //sfix24_En21
  parameter signed [23:0] coeff_b3_section5 = 24'b000010111111110111001010; //sfix24_En21
  parameter signed [23:0] coeff_a2_section5 = 24'b100000010110000101001001; //sfix24_En22
  parameter signed [23:0] coeff_a3_section5 = 24'b001111101111101101001010; //sfix24_En22
  parameter signed [23:0] coeff_b1_section6 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section6 = 24'b101010010001111011001110; //sfix24_En21
  parameter signed [23:0] coeff_b3_section6 = 24'b010011001000111000100001; //sfix24_En21
  parameter signed [23:0] coeff_a2_section6 = 24'b111001111000000110100100; //sfix24_En22
  parameter signed [23:0] coeff_a3_section6 = 24'b000001110110000100100111; //sfix24_En22
  parameter signed [23:0] coeff_b1_section7 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section7 = 24'b111001001000111101111110; //sfix24_En21
  parameter signed [23:0] coeff_b3_section7 = 24'b000100100100111010001001; //sfix24_En21
  parameter signed [23:0] coeff_a2_section7 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section7 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section8 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section8 = 24'b110011011010001000010010; //sfix24_En21
  parameter signed [23:0] coeff_b3_section8 = 24'b000100100101111111111011; //sfix24_En21
  parameter signed [23:0] coeff_a2_section8 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section8 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section9 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section9 = 24'b000010101110011010000111; //sfix24_En21
  parameter signed [23:0] coeff_b3_section9 = 24'b000000001001110001010100; //sfix24_En21
  parameter signed [23:0] coeff_a2_section9 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section9 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section10 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section10 = 24'b000010011011111111001111; //sfix24_En21
  parameter signed [23:0] coeff_b3_section10 = 24'b000000000001110110010111; //sfix24_En21
  parameter signed [23:0] coeff_a2_section10 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section10 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section11 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section11 = 24'b111111111011000011001001; //sfix24_En21
  parameter signed [23:0] coeff_b3_section11 = 24'b000000000000000110000100; //sfix24_En21
  parameter signed [23:0] coeff_a2_section11 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section11 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_b1_section12 = 24'b001000000000000000000000; //sfix24_En21
  parameter signed [23:0] coeff_b2_section12 = 24'b110111100110101100001000; //sfix24_En21
  parameter signed [23:0] coeff_b3_section12 = 24'b000000011001011001010100; //sfix24_En21
  parameter signed [23:0] coeff_a2_section12 = 24'b000000000000000000000000; //sfix24_En22
  parameter signed [23:0] coeff_a3_section12 = 24'b000000000000000000000000; //sfix24_En22
  // Signals
  reg  signed [23:0] input_register; // sfix24_En23
  wire signed [52:0] scale1; // sfix53_En57
  wire signed [47:0] mul_temp; // sfix48_En57
  wire signed [23:0] scaletypeconvert1; // sfix24_En28
  // Section 1 Signals 
  wire signed [39:0] a1sum1; // sfix40_En35
  wire signed [39:0] a2sum1; // sfix40_En35
  wire signed [39:0] b1sum1; // sfix40_En34
  wire signed [39:0] b2sum1; // sfix40_En34
  wire signed [23:0] typeconvert1; // sfix24_En23
  reg  signed [23:0] delay_section1 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv1; // sfix40_En35
  wire signed [47:0] a2mul1; // sfix48_En45
  wire signed [47:0] a3mul1; // sfix48_En45
  wire signed [47:0] b1mul1; // sfix48_En44
  wire signed [47:0] b2mul1; // sfix48_En44
  wire signed [47:0] b3mul1; // sfix48_En44
  wire signed [39:0] sub_cast; // sfix40_En35
  wire signed [39:0] sub_cast_1; // sfix40_En35
  wire signed [40:0] sub_temp; // sfix41_En35
  wire signed [39:0] sub_cast_2; // sfix40_En35
  wire signed [39:0] sub_cast_3; // sfix40_En35
  wire signed [40:0] sub_temp_1; // sfix41_En35
  wire signed [39:0] b1multypeconvert1; // sfix40_En34
  wire signed [39:0] add_cast; // sfix40_En34
  wire signed [39:0] add_cast_1; // sfix40_En34
  wire signed [40:0] add_temp; // sfix41_En34
  wire signed [39:0] add_cast_2; // sfix40_En34
  wire signed [39:0] add_cast_3; // sfix40_En34
  wire signed [40:0] add_temp_1; // sfix41_En34
  wire signed [39:0] section_result1; // sfix40_En35
  // Section 2 Signals 
  wire signed [39:0] a1sum2; // sfix40_En35
  wire signed [39:0] a2sum2; // sfix40_En35
  wire signed [39:0] b1sum2; // sfix40_En34
  wire signed [39:0] b2sum2; // sfix40_En34
  wire signed [23:0] typeconvert2; // sfix24_En23
  reg  signed [23:0] delay_section2 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv2; // sfix40_En35
  wire signed [47:0] a2mul2; // sfix48_En45
  wire signed [47:0] a3mul2; // sfix48_En45
  wire signed [47:0] b1mul2; // sfix48_En44
  wire signed [47:0] b2mul2; // sfix48_En44
  wire signed [47:0] b3mul2; // sfix48_En44
  wire signed [39:0] sub_cast_4; // sfix40_En35
  wire signed [39:0] sub_cast_5; // sfix40_En35
  wire signed [40:0] sub_temp_2; // sfix41_En35
  wire signed [39:0] sub_cast_6; // sfix40_En35
  wire signed [39:0] sub_cast_7; // sfix40_En35
  wire signed [40:0] sub_temp_3; // sfix41_En35
  wire signed [39:0] b1multypeconvert2; // sfix40_En34
  wire signed [39:0] add_cast_4; // sfix40_En34
  wire signed [39:0] add_cast_5; // sfix40_En34
  wire signed [40:0] add_temp_2; // sfix41_En34
  wire signed [39:0] add_cast_6; // sfix40_En34
  wire signed [39:0] add_cast_7; // sfix40_En34
  wire signed [40:0] add_temp_3; // sfix41_En34
  wire signed [39:0] section_result2; // sfix40_En35
  // Section 3 Signals 
  wire signed [39:0] a1sum3; // sfix40_En35
  wire signed [39:0] a2sum3; // sfix40_En35
  wire signed [39:0] b1sum3; // sfix40_En34
  wire signed [39:0] b2sum3; // sfix40_En34
  wire signed [23:0] typeconvert3; // sfix24_En23
  reg  signed [23:0] delay_section3 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv3; // sfix40_En35
  wire signed [47:0] a2mul3; // sfix48_En45
  wire signed [47:0] a3mul3; // sfix48_En45
  wire signed [47:0] b1mul3; // sfix48_En44
  wire signed [47:0] b2mul3; // sfix48_En44
  wire signed [47:0] b3mul3; // sfix48_En44
  wire signed [39:0] sub_cast_8; // sfix40_En35
  wire signed [39:0] sub_cast_9; // sfix40_En35
  wire signed [40:0] sub_temp_4; // sfix41_En35
  wire signed [39:0] sub_cast_10; // sfix40_En35
  wire signed [39:0] sub_cast_11; // sfix40_En35
  wire signed [40:0] sub_temp_5; // sfix41_En35
  wire signed [39:0] b1multypeconvert3; // sfix40_En34
  wire signed [39:0] add_cast_8; // sfix40_En34
  wire signed [39:0] add_cast_9; // sfix40_En34
  wire signed [40:0] add_temp_4; // sfix41_En34
  wire signed [39:0] add_cast_10; // sfix40_En34
  wire signed [39:0] add_cast_11; // sfix40_En34
  wire signed [40:0] add_temp_5; // sfix41_En34
  wire signed [39:0] section_result3; // sfix40_En35
  // Section 4 Signals 
  wire signed [39:0] a1sum4; // sfix40_En35
  wire signed [39:0] a2sum4; // sfix40_En35
  wire signed [39:0] b1sum4; // sfix40_En34
  wire signed [39:0] b2sum4; // sfix40_En34
  wire signed [23:0] typeconvert4; // sfix24_En23
  reg  signed [23:0] delay_section4 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv4; // sfix40_En35
  wire signed [47:0] a2mul4; // sfix48_En45
  wire signed [47:0] a3mul4; // sfix48_En45
  wire signed [47:0] b1mul4; // sfix48_En44
  wire signed [47:0] b2mul4; // sfix48_En44
  wire signed [47:0] b3mul4; // sfix48_En44
  wire signed [39:0] sub_cast_12; // sfix40_En35
  wire signed [39:0] sub_cast_13; // sfix40_En35
  wire signed [40:0] sub_temp_6; // sfix41_En35
  wire signed [39:0] sub_cast_14; // sfix40_En35
  wire signed [39:0] sub_cast_15; // sfix40_En35
  wire signed [40:0] sub_temp_7; // sfix41_En35
  wire signed [39:0] b1multypeconvert4; // sfix40_En34
  wire signed [39:0] add_cast_12; // sfix40_En34
  wire signed [39:0] add_cast_13; // sfix40_En34
  wire signed [40:0] add_temp_6; // sfix41_En34
  wire signed [39:0] add_cast_14; // sfix40_En34
  wire signed [39:0] add_cast_15; // sfix40_En34
  wire signed [40:0] add_temp_7; // sfix41_En34
  wire signed [39:0] section_result4; // sfix40_En35
  // Section 5 Signals 
  wire signed [39:0] a1sum5; // sfix40_En35
  wire signed [39:0] a2sum5; // sfix40_En35
  wire signed [39:0] b1sum5; // sfix40_En34
  wire signed [39:0] b2sum5; // sfix40_En34
  wire signed [23:0] typeconvert5; // sfix24_En23
  reg  signed [23:0] delay_section5 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv5; // sfix40_En35
  wire signed [47:0] a2mul5; // sfix48_En45
  wire signed [47:0] a3mul5; // sfix48_En45
  wire signed [47:0] b1mul5; // sfix48_En44
  wire signed [47:0] b2mul5; // sfix48_En44
  wire signed [47:0] b3mul5; // sfix48_En44
  wire signed [39:0] sub_cast_16; // sfix40_En35
  wire signed [39:0] sub_cast_17; // sfix40_En35
  wire signed [40:0] sub_temp_8; // sfix41_En35
  wire signed [39:0] sub_cast_18; // sfix40_En35
  wire signed [39:0] sub_cast_19; // sfix40_En35
  wire signed [40:0] sub_temp_9; // sfix41_En35
  wire signed [39:0] b1multypeconvert5; // sfix40_En34
  wire signed [39:0] add_cast_16; // sfix40_En34
  wire signed [39:0] add_cast_17; // sfix40_En34
  wire signed [40:0] add_temp_8; // sfix41_En34
  wire signed [39:0] add_cast_18; // sfix40_En34
  wire signed [39:0] add_cast_19; // sfix40_En34
  wire signed [40:0] add_temp_9; // sfix41_En34
  wire signed [39:0] section_result5; // sfix40_En35
  // Section 6 Signals 
  wire signed [39:0] a1sum6; // sfix40_En35
  wire signed [39:0] a2sum6; // sfix40_En35
  wire signed [39:0] b1sum6; // sfix40_En34
  wire signed [39:0] b2sum6; // sfix40_En34
  wire signed [23:0] typeconvert6; // sfix24_En23
  reg  signed [23:0] delay_section6 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv6; // sfix40_En35
  wire signed [47:0] a2mul6; // sfix48_En45
  wire signed [47:0] a3mul6; // sfix48_En45
  wire signed [47:0] b1mul6; // sfix48_En44
  wire signed [47:0] b2mul6; // sfix48_En44
  wire signed [47:0] b3mul6; // sfix48_En44
  wire signed [39:0] sub_cast_20; // sfix40_En35
  wire signed [39:0] sub_cast_21; // sfix40_En35
  wire signed [40:0] sub_temp_10; // sfix41_En35
  wire signed [39:0] sub_cast_22; // sfix40_En35
  wire signed [39:0] sub_cast_23; // sfix40_En35
  wire signed [40:0] sub_temp_11; // sfix41_En35
  wire signed [39:0] b1multypeconvert6; // sfix40_En34
  wire signed [39:0] add_cast_20; // sfix40_En34
  wire signed [39:0] add_cast_21; // sfix40_En34
  wire signed [40:0] add_temp_10; // sfix41_En34
  wire signed [39:0] add_cast_22; // sfix40_En34
  wire signed [39:0] add_cast_23; // sfix40_En34
  wire signed [40:0] add_temp_11; // sfix41_En34
  wire signed [39:0] section_result6; // sfix40_En35
  // Section 7 Signals 
  wire signed [39:0] a1sum7; // sfix40_En35
  wire signed [39:0] b1sum7; // sfix40_En34
  wire signed [39:0] b2sum7; // sfix40_En34
  wire signed [23:0] typeconvert7; // sfix24_En23
  reg  signed [23:0] delay_section7 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv7; // sfix40_En35
  wire signed [47:0] b1mul7; // sfix48_En44
  wire signed [47:0] b2mul7; // sfix48_En44
  wire signed [47:0] b3mul7; // sfix48_En44
  wire signed [39:0] b1multypeconvert7; // sfix40_En34
  wire signed [39:0] add_cast_24; // sfix40_En34
  wire signed [39:0] add_cast_25; // sfix40_En34
  wire signed [40:0] add_temp_12; // sfix41_En34
  wire signed [39:0] add_cast_26; // sfix40_En34
  wire signed [39:0] add_cast_27; // sfix40_En34
  wire signed [40:0] add_temp_13; // sfix41_En34
  wire signed [39:0] section_result7; // sfix40_En35
  // Section 8 Signals 
  wire signed [39:0] a1sum8; // sfix40_En35
  wire signed [39:0] b1sum8; // sfix40_En34
  wire signed [39:0] b2sum8; // sfix40_En34
  wire signed [23:0] typeconvert8; // sfix24_En23
  reg  signed [23:0] delay_section8 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv8; // sfix40_En35
  wire signed [47:0] b1mul8; // sfix48_En44
  wire signed [47:0] b2mul8; // sfix48_En44
  wire signed [47:0] b3mul8; // sfix48_En44
  wire signed [39:0] b1multypeconvert8; // sfix40_En34
  wire signed [39:0] add_cast_28; // sfix40_En34
  wire signed [39:0] add_cast_29; // sfix40_En34
  wire signed [40:0] add_temp_14; // sfix41_En34
  wire signed [39:0] add_cast_30; // sfix40_En34
  wire signed [39:0] add_cast_31; // sfix40_En34
  wire signed [40:0] add_temp_15; // sfix41_En34
  wire signed [39:0] section_result8; // sfix40_En35
  // Section 9 Signals 
  wire signed [39:0] a1sum9; // sfix40_En35
  wire signed [39:0] b1sum9; // sfix40_En34
  wire signed [39:0] b2sum9; // sfix40_En34
  wire signed [23:0] typeconvert9; // sfix24_En23
  reg  signed [23:0] delay_section9 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv9; // sfix40_En35
  wire signed [47:0] b1mul9; // sfix48_En44
  wire signed [47:0] b2mul9; // sfix48_En44
  wire signed [47:0] b3mul9; // sfix48_En44
  wire signed [39:0] b1multypeconvert9; // sfix40_En34
  wire signed [39:0] add_cast_32; // sfix40_En34
  wire signed [39:0] add_cast_33; // sfix40_En34
  wire signed [40:0] add_temp_16; // sfix41_En34
  wire signed [39:0] add_cast_34; // sfix40_En34
  wire signed [39:0] add_cast_35; // sfix40_En34
  wire signed [40:0] add_temp_17; // sfix41_En34
  wire signed [39:0] section_result9; // sfix40_En35
  // Section 10 Signals 
  wire signed [39:0] a1sum10; // sfix40_En35
  wire signed [39:0] b1sum10; // sfix40_En34
  wire signed [39:0] b2sum10; // sfix40_En34
  wire signed [23:0] typeconvert10; // sfix24_En23
  reg  signed [23:0] delay_section10 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv10; // sfix40_En35
  wire signed [47:0] b1mul10; // sfix48_En44
  wire signed [47:0] b2mul10; // sfix48_En44
  wire signed [47:0] b3mul10; // sfix48_En44
  wire signed [39:0] b1multypeconvert10; // sfix40_En34
  wire signed [39:0] add_cast_36; // sfix40_En34
  wire signed [39:0] add_cast_37; // sfix40_En34
  wire signed [40:0] add_temp_18; // sfix41_En34
  wire signed [39:0] add_cast_38; // sfix40_En34
  wire signed [39:0] add_cast_39; // sfix40_En34
  wire signed [40:0] add_temp_19; // sfix41_En34
  wire signed [39:0] section_result10; // sfix40_En35
  // Section 11 Signals 
  wire signed [39:0] a1sum11; // sfix40_En35
  wire signed [39:0] b1sum11; // sfix40_En34
  wire signed [39:0] b2sum11; // sfix40_En34
  wire signed [23:0] typeconvert11; // sfix24_En23
  reg  signed [23:0] delay_section11 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv11; // sfix40_En35
  wire signed [47:0] b1mul11; // sfix48_En44
  wire signed [47:0] b2mul11; // sfix48_En44
  wire signed [47:0] b3mul11; // sfix48_En44
  wire signed [39:0] b1multypeconvert11; // sfix40_En34
  wire signed [39:0] add_cast_40; // sfix40_En34
  wire signed [39:0] add_cast_41; // sfix40_En34
  wire signed [40:0] add_temp_20; // sfix41_En34
  wire signed [39:0] add_cast_42; // sfix40_En34
  wire signed [39:0] add_cast_43; // sfix40_En34
  wire signed [40:0] add_temp_21; // sfix41_En34
  wire signed [39:0] section_result11; // sfix40_En35
  // Section 12 Signals 
  wire signed [39:0] a1sum12; // sfix40_En35
  wire signed [39:0] b1sum12; // sfix40_En34
  wire signed [39:0] b2sum12; // sfix40_En34
  wire signed [23:0] typeconvert12; // sfix24_En23
  reg  signed [23:0] delay_section12 [0:1] ; // sfix24_En23
  wire signed [39:0] inputconv12; // sfix40_En35
  wire signed [47:0] b1mul12; // sfix48_En44
  wire signed [47:0] b2mul12; // sfix48_En44
  wire signed [47:0] b3mul12; // sfix48_En44
  wire signed [39:0] b1multypeconvert12; // sfix40_En34
  wire signed [39:0] add_cast_44; // sfix40_En34
  wire signed [39:0] add_cast_45; // sfix40_En34
  wire signed [40:0] add_temp_22; // sfix41_En34
  wire signed [39:0] add_cast_46; // sfix40_En34
  wire signed [39:0] add_cast_47; // sfix40_En34
  wire signed [40:0] add_temp_23; // sfix41_En34
  wire signed [23:0] output_typeconvert; // sfix24_En18
  reg  signed [23:0] output_register; // sfix24_En18

  // Block Statements
  always @ (posedge clk or posedge reset)
    begin: input_reg_process
      if (reset == 1'b1) begin
        input_register <= 0;
      end
      else begin
        if (clk_enable == 1'b1) begin
          input_register <= filter_in;
        end
      end
    end // input_reg_process

  assign mul_temp = input_register * scaleconst1;
  assign scale1 = $signed({{5{mul_temp[47]}}, mul_temp});

  assign scaletypeconvert1 = (scale1[52:0] + {scale1[29], {28{~scale1[29]}}})>>>29;

  //   ------------------ Section 1 ------------------

  assign typeconvert1 = (a1sum1[35:0] + {a1sum1[12], {11{~a1sum1[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section1
      if (reset == 1'b1) begin
        delay_section1[0] <= 24'b000000000000000000000000;
        delay_section1[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section1[1] <= delay_section1[0];
          delay_section1[0] <= typeconvert1;
        end
      end
    end // delay_process_section1

  assign inputconv1 = $signed({scaletypeconvert1[23:0], 7'b0000000});

  assign a2mul1 = delay_section1[0] * coeff_a2_section1;

  assign a3mul1 = delay_section1[1] * coeff_a3_section1;

  assign b1mul1 = $signed({typeconvert1[23:0], 21'b000000000000000000000});

  assign b2mul1 = delay_section1[0] * coeff_b2_section1;

  assign b3mul1 = delay_section1[1] * coeff_b3_section1;

  assign sub_cast = inputconv1;
  assign sub_cast_1 = ({{2{a2mul1[47]}}, a2mul1[47:0]} + {a2mul1[10], {9{~a2mul1[10]}}})>>>10;
  assign sub_temp = sub_cast - sub_cast_1;
  assign a2sum1 = sub_temp[39:0];

  assign sub_cast_2 = a2sum1;
  assign sub_cast_3 = ({{2{a3mul1[47]}}, a3mul1[47:0]} + {a3mul1[10], {9{~a3mul1[10]}}})>>>10;
  assign sub_temp_1 = sub_cast_2 - sub_cast_3;
  assign a1sum1 = sub_temp_1[39:0];

  assign b1multypeconvert1 = ({{2{b1mul1[47]}}, b1mul1[47:0]} + {b1mul1[10], {9{~b1mul1[10]}}})>>>10;

  assign add_cast = b1multypeconvert1;
  assign add_cast_1 = ({{2{b2mul1[47]}}, b2mul1[47:0]} + {b2mul1[10], {9{~b2mul1[10]}}})>>>10;
  assign add_temp = add_cast + add_cast_1;
  assign b2sum1 = add_temp[39:0];

  assign add_cast_2 = b2sum1;
  assign add_cast_3 = ({{2{b3mul1[47]}}, b3mul1[47:0]} + {b3mul1[10], {9{~b3mul1[10]}}})>>>10;
  assign add_temp_1 = add_cast_2 + add_cast_3;
  assign b1sum1 = add_temp_1[39:0];

  assign section_result1 = $signed({b1sum1[38:0], 1'b0});

  //   ------------------ Section 2 ------------------

  assign typeconvert2 = (a1sum2[35:0] + {a1sum2[12], {11{~a1sum2[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section2
      if (reset == 1'b1) begin
        delay_section2[0] <= 24'b000000000000000000000000;
        delay_section2[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section2[1] <= delay_section2[0];
          delay_section2[0] <= typeconvert2;
        end
      end
    end // delay_process_section2

  assign inputconv2 = section_result1;

  assign a2mul2 = delay_section2[0] * coeff_a2_section2;

  assign a3mul2 = delay_section2[1] * coeff_a3_section2;

  assign b1mul2 = $signed({typeconvert2[23:0], 21'b000000000000000000000});

  assign b2mul2 = delay_section2[0] * coeff_b2_section2;

  assign b3mul2 = delay_section2[1] * coeff_b3_section2;

  assign sub_cast_4 = inputconv2;
  assign sub_cast_5 = ({{2{a2mul2[47]}}, a2mul2[47:0]} + {a2mul2[10], {9{~a2mul2[10]}}})>>>10;
  assign sub_temp_2 = sub_cast_4 - sub_cast_5;
  assign a2sum2 = sub_temp_2[39:0];

  assign sub_cast_6 = a2sum2;
  assign sub_cast_7 = ({{2{a3mul2[47]}}, a3mul2[47:0]} + {a3mul2[10], {9{~a3mul2[10]}}})>>>10;
  assign sub_temp_3 = sub_cast_6 - sub_cast_7;
  assign a1sum2 = sub_temp_3[39:0];

  assign b1multypeconvert2 = ({{2{b1mul2[47]}}, b1mul2[47:0]} + {b1mul2[10], {9{~b1mul2[10]}}})>>>10;

  assign add_cast_4 = b1multypeconvert2;
  assign add_cast_5 = ({{2{b2mul2[47]}}, b2mul2[47:0]} + {b2mul2[10], {9{~b2mul2[10]}}})>>>10;
  assign add_temp_2 = add_cast_4 + add_cast_5;
  assign b2sum2 = add_temp_2[39:0];

  assign add_cast_6 = b2sum2;
  assign add_cast_7 = ({{2{b3mul2[47]}}, b3mul2[47:0]} + {b3mul2[10], {9{~b3mul2[10]}}})>>>10;
  assign add_temp_3 = add_cast_6 + add_cast_7;
  assign b1sum2 = add_temp_3[39:0];

  assign section_result2 = $signed({b1sum2[38:0], 1'b0});

  //   ------------------ Section 3 ------------------

  assign typeconvert3 = (a1sum3[35:0] + {a1sum3[12], {11{~a1sum3[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section3
      if (reset == 1'b1) begin
        delay_section3[0] <= 24'b000000000000000000000000;
        delay_section3[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section3[1] <= delay_section3[0];
          delay_section3[0] <= typeconvert3;
        end
      end
    end // delay_process_section3

  assign inputconv3 = section_result2;

  assign a2mul3 = delay_section3[0] * coeff_a2_section3;

  assign a3mul3 = delay_section3[1] * coeff_a3_section3;

  assign b1mul3 = $signed({typeconvert3[23:0], 21'b000000000000000000000});

  assign b2mul3 = delay_section3[0] * coeff_b2_section3;

  assign b3mul3 = delay_section3[1] * coeff_b3_section3;

  assign sub_cast_8 = inputconv3;
  assign sub_cast_9 = ({{2{a2mul3[47]}}, a2mul3[47:0]} + {a2mul3[10], {9{~a2mul3[10]}}})>>>10;
  assign sub_temp_4 = sub_cast_8 - sub_cast_9;
  assign a2sum3 = sub_temp_4[39:0];

  assign sub_cast_10 = a2sum3;
  assign sub_cast_11 = ({{2{a3mul3[47]}}, a3mul3[47:0]} + {a3mul3[10], {9{~a3mul3[10]}}})>>>10;
  assign sub_temp_5 = sub_cast_10 - sub_cast_11;
  assign a1sum3 = sub_temp_5[39:0];

  assign b1multypeconvert3 = ({{2{b1mul3[47]}}, b1mul3[47:0]} + {b1mul3[10], {9{~b1mul3[10]}}})>>>10;

  assign add_cast_8 = b1multypeconvert3;
  assign add_cast_9 = ({{2{b2mul3[47]}}, b2mul3[47:0]} + {b2mul3[10], {9{~b2mul3[10]}}})>>>10;
  assign add_temp_4 = add_cast_8 + add_cast_9;
  assign b2sum3 = add_temp_4[39:0];

  assign add_cast_10 = b2sum3;
  assign add_cast_11 = ({{2{b3mul3[47]}}, b3mul3[47:0]} + {b3mul3[10], {9{~b3mul3[10]}}})>>>10;
  assign add_temp_5 = add_cast_10 + add_cast_11;
  assign b1sum3 = add_temp_5[39:0];

  assign section_result3 = $signed({b1sum3[38:0], 1'b0});

  //   ------------------ Section 4 ------------------

  assign typeconvert4 = (a1sum4[35:0] + {a1sum4[12], {11{~a1sum4[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section4
      if (reset == 1'b1) begin
        delay_section4[0] <= 24'b000000000000000000000000;
        delay_section4[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section4[1] <= delay_section4[0];
          delay_section4[0] <= typeconvert4;
        end
      end
    end // delay_process_section4

  assign inputconv4 = section_result3;

  assign a2mul4 = delay_section4[0] * coeff_a2_section4;

  assign a3mul4 = delay_section4[1] * coeff_a3_section4;

  assign b1mul4 = $signed({typeconvert4[23:0], 21'b000000000000000000000});

  assign b2mul4 = delay_section4[0] * coeff_b2_section4;

  assign b3mul4 = delay_section4[1] * coeff_b3_section4;

  assign sub_cast_12 = inputconv4;
  assign sub_cast_13 = ({{2{a2mul4[47]}}, a2mul4[47:0]} + {a2mul4[10], {9{~a2mul4[10]}}})>>>10;
  assign sub_temp_6 = sub_cast_12 - sub_cast_13;
  assign a2sum4 = sub_temp_6[39:0];

  assign sub_cast_14 = a2sum4;
  assign sub_cast_15 = ({{2{a3mul4[47]}}, a3mul4[47:0]} + {a3mul4[10], {9{~a3mul4[10]}}})>>>10;
  assign sub_temp_7 = sub_cast_14 - sub_cast_15;
  assign a1sum4 = sub_temp_7[39:0];

  assign b1multypeconvert4 = ({{2{b1mul4[47]}}, b1mul4[47:0]} + {b1mul4[10], {9{~b1mul4[10]}}})>>>10;

  assign add_cast_12 = b1multypeconvert4;
  assign add_cast_13 = ({{2{b2mul4[47]}}, b2mul4[47:0]} + {b2mul4[10], {9{~b2mul4[10]}}})>>>10;
  assign add_temp_6 = add_cast_12 + add_cast_13;
  assign b2sum4 = add_temp_6[39:0];

  assign add_cast_14 = b2sum4;
  assign add_cast_15 = ({{2{b3mul4[47]}}, b3mul4[47:0]} + {b3mul4[10], {9{~b3mul4[10]}}})>>>10;
  assign add_temp_7 = add_cast_14 + add_cast_15;
  assign b1sum4 = add_temp_7[39:0];

  assign section_result4 = $signed({b1sum4[38:0], 1'b0});

  //   ------------------ Section 5 ------------------

  assign typeconvert5 = (a1sum5[35:0] + {a1sum5[12], {11{~a1sum5[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section5
      if (reset == 1'b1) begin
        delay_section5[0] <= 24'b000000000000000000000000;
        delay_section5[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section5[1] <= delay_section5[0];
          delay_section5[0] <= typeconvert5;
        end
      end
    end // delay_process_section5

  assign inputconv5 = section_result4;

  assign a2mul5 = delay_section5[0] * coeff_a2_section5;

  assign a3mul5 = delay_section5[1] * coeff_a3_section5;

  assign b1mul5 = $signed({typeconvert5[23:0], 21'b000000000000000000000});

  assign b2mul5 = delay_section5[0] * coeff_b2_section5;

  assign b3mul5 = delay_section5[1] * coeff_b3_section5;

  assign sub_cast_16 = inputconv5;
  assign sub_cast_17 = ({{2{a2mul5[47]}}, a2mul5[47:0]} + {a2mul5[10], {9{~a2mul5[10]}}})>>>10;
  assign sub_temp_8 = sub_cast_16 - sub_cast_17;
  assign a2sum5 = sub_temp_8[39:0];

  assign sub_cast_18 = a2sum5;
  assign sub_cast_19 = ({{2{a3mul5[47]}}, a3mul5[47:0]} + {a3mul5[10], {9{~a3mul5[10]}}})>>>10;
  assign sub_temp_9 = sub_cast_18 - sub_cast_19;
  assign a1sum5 = sub_temp_9[39:0];

  assign b1multypeconvert5 = ({{2{b1mul5[47]}}, b1mul5[47:0]} + {b1mul5[10], {9{~b1mul5[10]}}})>>>10;

  assign add_cast_16 = b1multypeconvert5;
  assign add_cast_17 = ({{2{b2mul5[47]}}, b2mul5[47:0]} + {b2mul5[10], {9{~b2mul5[10]}}})>>>10;
  assign add_temp_8 = add_cast_16 + add_cast_17;
  assign b2sum5 = add_temp_8[39:0];

  assign add_cast_18 = b2sum5;
  assign add_cast_19 = ({{2{b3mul5[47]}}, b3mul5[47:0]} + {b3mul5[10], {9{~b3mul5[10]}}})>>>10;
  assign add_temp_9 = add_cast_18 + add_cast_19;
  assign b1sum5 = add_temp_9[39:0];

  assign section_result5 = $signed({b1sum5[38:0], 1'b0});

  //   ------------------ Section 6 ------------------

  assign typeconvert6 = (a1sum6[35:0] + {a1sum6[12], {11{~a1sum6[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section6
      if (reset == 1'b1) begin
        delay_section6[0] <= 24'b000000000000000000000000;
        delay_section6[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section6[1] <= delay_section6[0];
          delay_section6[0] <= typeconvert6;
        end
      end
    end // delay_process_section6

  assign inputconv6 = section_result5;

  assign a2mul6 = delay_section6[0] * coeff_a2_section6;

  assign a3mul6 = delay_section6[1] * coeff_a3_section6;

  assign b1mul6 = $signed({typeconvert6[23:0], 21'b000000000000000000000});

  assign b2mul6 = delay_section6[0] * coeff_b2_section6;

  assign b3mul6 = delay_section6[1] * coeff_b3_section6;

  assign sub_cast_20 = inputconv6;
  assign sub_cast_21 = ({{2{a2mul6[47]}}, a2mul6[47:0]} + {a2mul6[10], {9{~a2mul6[10]}}})>>>10;
  assign sub_temp_10 = sub_cast_20 - sub_cast_21;
  assign a2sum6 = sub_temp_10[39:0];

  assign sub_cast_22 = a2sum6;
  assign sub_cast_23 = ({{2{a3mul6[47]}}, a3mul6[47:0]} + {a3mul6[10], {9{~a3mul6[10]}}})>>>10;
  assign sub_temp_11 = sub_cast_22 - sub_cast_23;
  assign a1sum6 = sub_temp_11[39:0];

  assign b1multypeconvert6 = ({{2{b1mul6[47]}}, b1mul6[47:0]} + {b1mul6[10], {9{~b1mul6[10]}}})>>>10;

  assign add_cast_20 = b1multypeconvert6;
  assign add_cast_21 = ({{2{b2mul6[47]}}, b2mul6[47:0]} + {b2mul6[10], {9{~b2mul6[10]}}})>>>10;
  assign add_temp_10 = add_cast_20 + add_cast_21;
  assign b2sum6 = add_temp_10[39:0];

  assign add_cast_22 = b2sum6;
  assign add_cast_23 = ({{2{b3mul6[47]}}, b3mul6[47:0]} + {b3mul6[10], {9{~b3mul6[10]}}})>>>10;
  assign add_temp_11 = add_cast_22 + add_cast_23;
  assign b1sum6 = add_temp_11[39:0];

  assign section_result6 = $signed({b1sum6[38:0], 1'b0});

  //   ------------------ Section 7 ------------------

  assign typeconvert7 = (a1sum7[35:0] + {a1sum7[12], {11{~a1sum7[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section7
      if (reset == 1'b1) begin
        delay_section7[0] <= 24'b000000000000000000000000;
        delay_section7[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section7[1] <= delay_section7[0];
          delay_section7[0] <= typeconvert7;
        end
      end
    end // delay_process_section7

  assign inputconv7 = section_result6;

  assign b1mul7 = $signed({typeconvert7[23:0], 21'b000000000000000000000});

  assign b2mul7 = delay_section7[0] * coeff_b2_section7;

  assign b3mul7 = delay_section7[1] * coeff_b3_section7;

  assign a1sum7 = inputconv7;

  assign b1multypeconvert7 = ({{2{b1mul7[47]}}, b1mul7[47:0]} + {b1mul7[10], {9{~b1mul7[10]}}})>>>10;

  assign add_cast_24 = b1multypeconvert7;
  assign add_cast_25 = ({{2{b2mul7[47]}}, b2mul7[47:0]} + {b2mul7[10], {9{~b2mul7[10]}}})>>>10;
  assign add_temp_12 = add_cast_24 + add_cast_25;
  assign b2sum7 = add_temp_12[39:0];

  assign add_cast_26 = b2sum7;
  assign add_cast_27 = ({{2{b3mul7[47]}}, b3mul7[47:0]} + {b3mul7[10], {9{~b3mul7[10]}}})>>>10;
  assign add_temp_13 = add_cast_26 + add_cast_27;
  assign b1sum7 = add_temp_13[39:0];

  assign section_result7 = $signed({b1sum7[38:0], 1'b0});

  //   ------------------ Section 8 ------------------

  assign typeconvert8 = (a1sum8[35:0] + {a1sum8[12], {11{~a1sum8[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section8
      if (reset == 1'b1) begin
        delay_section8[0] <= 24'b000000000000000000000000;
        delay_section8[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section8[1] <= delay_section8[0];
          delay_section8[0] <= typeconvert8;
        end
      end
    end // delay_process_section8

  assign inputconv8 = section_result7;

  assign b1mul8 = $signed({typeconvert8[23:0], 21'b000000000000000000000});

  assign b2mul8 = delay_section8[0] * coeff_b2_section8;

  assign b3mul8 = delay_section8[1] * coeff_b3_section8;

  assign a1sum8 = inputconv8;

  assign b1multypeconvert8 = ({{2{b1mul8[47]}}, b1mul8[47:0]} + {b1mul8[10], {9{~b1mul8[10]}}})>>>10;

  assign add_cast_28 = b1multypeconvert8;
  assign add_cast_29 = ({{2{b2mul8[47]}}, b2mul8[47:0]} + {b2mul8[10], {9{~b2mul8[10]}}})>>>10;
  assign add_temp_14 = add_cast_28 + add_cast_29;
  assign b2sum8 = add_temp_14[39:0];

  assign add_cast_30 = b2sum8;
  assign add_cast_31 = ({{2{b3mul8[47]}}, b3mul8[47:0]} + {b3mul8[10], {9{~b3mul8[10]}}})>>>10;
  assign add_temp_15 = add_cast_30 + add_cast_31;
  assign b1sum8 = add_temp_15[39:0];

  assign section_result8 = $signed({b1sum8[38:0], 1'b0});

  //   ------------------ Section 9 ------------------

  assign typeconvert9 = (a1sum9[35:0] + {a1sum9[12], {11{~a1sum9[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section9
      if (reset == 1'b1) begin
        delay_section9[0] <= 24'b000000000000000000000000;
        delay_section9[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section9[1] <= delay_section9[0];
          delay_section9[0] <= typeconvert9;
        end
      end
    end // delay_process_section9

  assign inputconv9 = section_result8;

  assign b1mul9 = $signed({typeconvert9[23:0], 21'b000000000000000000000});

  assign b2mul9 = delay_section9[0] * coeff_b2_section9;

  assign b3mul9 = delay_section9[1] * coeff_b3_section9;

  assign a1sum9 = inputconv9;

  assign b1multypeconvert9 = ({{2{b1mul9[47]}}, b1mul9[47:0]} + {b1mul9[10], {9{~b1mul9[10]}}})>>>10;

  assign add_cast_32 = b1multypeconvert9;
  assign add_cast_33 = ({{2{b2mul9[47]}}, b2mul9[47:0]} + {b2mul9[10], {9{~b2mul9[10]}}})>>>10;
  assign add_temp_16 = add_cast_32 + add_cast_33;
  assign b2sum9 = add_temp_16[39:0];

  assign add_cast_34 = b2sum9;
  assign add_cast_35 = ({{2{b3mul9[47]}}, b3mul9[47:0]} + {b3mul9[10], {9{~b3mul9[10]}}})>>>10;
  assign add_temp_17 = add_cast_34 + add_cast_35;
  assign b1sum9 = add_temp_17[39:0];

  assign section_result9 = $signed({b1sum9[38:0], 1'b0});

  //   ------------------ Section 10 ------------------

  assign typeconvert10 = (a1sum10[35:0] + {a1sum10[12], {11{~a1sum10[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section10
      if (reset == 1'b1) begin
        delay_section10[0] <= 24'b000000000000000000000000;
        delay_section10[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section10[1] <= delay_section10[0];
          delay_section10[0] <= typeconvert10;
        end
      end
    end // delay_process_section10

  assign inputconv10 = section_result9;

  assign b1mul10 = $signed({typeconvert10[23:0], 21'b000000000000000000000});

  assign b2mul10 = delay_section10[0] * coeff_b2_section10;

  assign b3mul10 = delay_section10[1] * coeff_b3_section10;

  assign a1sum10 = inputconv10;

  assign b1multypeconvert10 = ({{2{b1mul10[47]}}, b1mul10[47:0]} + {b1mul10[10], {9{~b1mul10[10]}}})>>>10;

  assign add_cast_36 = b1multypeconvert10;
  assign add_cast_37 = ({{2{b2mul10[47]}}, b2mul10[47:0]} + {b2mul10[10], {9{~b2mul10[10]}}})>>>10;
  assign add_temp_18 = add_cast_36 + add_cast_37;
  assign b2sum10 = add_temp_18[39:0];

  assign add_cast_38 = b2sum10;
  assign add_cast_39 = ({{2{b3mul10[47]}}, b3mul10[47:0]} + {b3mul10[10], {9{~b3mul10[10]}}})>>>10;
  assign add_temp_19 = add_cast_38 + add_cast_39;
  assign b1sum10 = add_temp_19[39:0];

  assign section_result10 = $signed({b1sum10[38:0], 1'b0});

  //   ------------------ Section 11 ------------------

  assign typeconvert11 = (a1sum11[35:0] + {a1sum11[12], {11{~a1sum11[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section11
      if (reset == 1'b1) begin
        delay_section11[0] <= 24'b000000000000000000000000;
        delay_section11[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section11[1] <= delay_section11[0];
          delay_section11[0] <= typeconvert11;
        end
      end
    end // delay_process_section11

  assign inputconv11 = section_result10;

  assign b1mul11 = $signed({typeconvert11[23:0], 21'b000000000000000000000});

  assign b2mul11 = delay_section11[0] * coeff_b2_section11;

  assign b3mul11 = delay_section11[1] * coeff_b3_section11;

  assign a1sum11 = inputconv11;

  assign b1multypeconvert11 = ({{2{b1mul11[47]}}, b1mul11[47:0]} + {b1mul11[10], {9{~b1mul11[10]}}})>>>10;

  assign add_cast_40 = b1multypeconvert11;
  assign add_cast_41 = ({{2{b2mul11[47]}}, b2mul11[47:0]} + {b2mul11[10], {9{~b2mul11[10]}}})>>>10;
  assign add_temp_20 = add_cast_40 + add_cast_41;
  assign b2sum11 = add_temp_20[39:0];

  assign add_cast_42 = b2sum11;
  assign add_cast_43 = ({{2{b3mul11[47]}}, b3mul11[47:0]} + {b3mul11[10], {9{~b3mul11[10]}}})>>>10;
  assign add_temp_21 = add_cast_42 + add_cast_43;
  assign b1sum11 = add_temp_21[39:0];

  assign section_result11 = $signed({b1sum11[38:0], 1'b0});

  //   ------------------ Section 12 ------------------

  assign typeconvert12 = (a1sum12[35:0] + {a1sum12[12], {11{~a1sum12[12]}}})>>>12;

  always @ (posedge clk or posedge reset)
    begin: delay_process_section12
      if (reset == 1'b1) begin
        delay_section12[0] <= 24'b000000000000000000000000;
        delay_section12[1] <= 24'b000000000000000000000000;
      end
      else begin
        if (clk_enable == 1'b1) begin
          delay_section12[1] <= delay_section12[0];
          delay_section12[0] <= typeconvert12;
        end
      end
    end // delay_process_section12

  assign inputconv12 = section_result11;

  assign b1mul12 = $signed({typeconvert12[23:0], 21'b000000000000000000000});

  assign b2mul12 = delay_section12[0] * coeff_b2_section12;

  assign b3mul12 = delay_section12[1] * coeff_b3_section12;

  assign a1sum12 = inputconv12;

  assign b1multypeconvert12 = ({{2{b1mul12[47]}}, b1mul12[47:0]} + {b1mul12[10], {9{~b1mul12[10]}}})>>>10;

  assign add_cast_44 = b1multypeconvert12;
  assign add_cast_45 = ({{2{b2mul12[47]}}, b2mul12[47:0]} + {b2mul12[10], {9{~b2mul12[10]}}})>>>10;
  assign add_temp_22 = add_cast_44 + add_cast_45;
  assign b2sum12 = add_temp_22[39:0];

  assign add_cast_46 = b2sum12;
  assign add_cast_47 = ({{2{b3mul12[47]}}, b3mul12[47:0]} + {b3mul12[10], {9{~b3mul12[10]}}})>>>10;
  assign add_temp_23 = add_cast_46 + add_cast_47;
  assign b1sum12 = add_temp_23[39:0];

  assign output_typeconvert = (b1sum12[39:0] + {b1sum12[16], {15{~b1sum12[16]}}})>>>16;

  always @ (posedge clk or posedge reset)
    begin: Output_Register_process
      if (reset == 1'b1) begin
        output_register <= 0;
      end
      else begin
        if (clk_enable == 1'b1) begin
          output_register <= output_typeconvert;
        end
      end
    end // Output_Register_process

  // Assignment Statements
  assign filter_out = output_register;
endmodule  // bandpass_leastPth_ver

module MidiProcessor(
	input CLOCK_50,
	input MIDI_RX,
	output reg isNoteOn,
	output reg [23:0] noteSampleTicks,
	output reg [7:0] modulationValue
);

reg [3:0] status = 0;
reg [3:0] channel = 0;
reg [7:0] dataByte0 = 0;
reg [7:0] dataByte1 = 0;
reg [7:0] dataByte2 = 0;
reg [7:0] dataBytesReceivedCount = 0;
reg isDataByteAvailable = 0;
reg [7:0] midiNoteNumber = 0;
reg [7:0] controllerNumber = 0;

wire isByteAvailable;
wire [7:0] byteValue;
wire [23:0] sampleTicks;

//MidiByteReader midiByteReader(CLOCK_50, MIDI_RX, isByteAvailable, byteValue);
//MidiNoteNumberToSampleTicks midiNoteNumberToSampleTicks(midiNoteNumber, sampleTicks);

always @(posedge CLOCK_50)
begin
	if (isByteAvailable == 1'b1)
		begin
			if (byteValue < 8'h80)  // Data byte
				begin
					case (dataBytesReceivedCount)
						0:
							begin
								dataByte0 <= byteValue;
								dataBytesReceivedCount <= 8'd1;
								isDataByteAvailable <= 1'b1;
							end
						1:
							begin
								dataByte1 <= byteValue;
								dataBytesReceivedCount <= 8'd2;
								isDataByteAvailable <= 1'b1;
							end
						2:
							begin
								dataByte2 <= byteValue;
								dataBytesReceivedCount <= 8'd3;
								isDataByteAvailable <= 1'b1;
							end
					endcase
				end
			else  // Status byte
				begin
					status <= byteValue[7:4];
					channel <= byteValue[3:0];
					dataBytesReceivedCount <= 0;
				end
		end
	else if (isDataByteAvailable == 1'b1)
		begin
			isDataByteAvailable <= 1'b0;
		
			case (status)
				4'h8:  // Note Off
					if (dataBytesReceivedCount == 2)
						begin
							if (midiNoteNumber == dataByte0)
								begin
									dataBytesReceivedCount <= 0;
									isNoteOn <= 1'b0;
								end
						end
				4'h9:  // Note On
					case (dataBytesReceivedCount)
						1:
							midiNoteNumber <= dataByte0;
						2:
							begin
								dataBytesReceivedCount <= 0;

								if (dataByte1 == 0)
									begin
										// Zero velocity is like Note Off
										isNoteOn <= 1'b0;										
									end
								else
									begin
										isNoteOn <= 1'b1;
										noteSampleTicks <= sampleTicks;
									end
							end
					endcase
				4'hB:  // Controller Change
					case (dataBytesReceivedCount)
						1:
							controllerNumber <= dataByte0;
						2:
							begin
								if (controllerNumber == 8'd1)
									begin
										dataBytesReceivedCount <= 0;
										modulationValue <= dataByte1;
									end
							end
					endcase
			endcase
		end
end

endmodule

module Synthesizer(
	input CLOCK_50,
	input isNoteOn,
	input [23:0] noteSampleTicks,
	input [7:0] modulationValue,
	output reg i2sBitClock,
	output reg i2sSoundData,
	output reg i2sLeftRightSelect
);

// 50,000,000 / 44,100 / 16 / 2 / 2 (DE0 Nano clock / sample rate / bits per sample / channels / edges);
localparam i2sTicks = 8'd18;  // 17.7154195

reg [11:0] i2sCount = 0;
reg [23:0] noteSampleCount = 0;
reg [7:0] bitCount = 15;
reg [7:0] sampleIndex = 0;
reg [7:0] waveTableIndex = 0;
reg [7:0] modulation = 0;
reg isSamplePlaying = 0;
reg isSoundPlaying = 0;

wire [15:0] waveTableSample0;
wire [15:0] waveTableSample1;
wire [15:0] waveTableSample2;
wire [15:0] renderedSample;

//WaveTable0Rom waveTable0Rom(waveTableIndex, CLOCK_50, waveTableSample0);
//WaveTable1Rom waveTable1Rom(waveTableIndex, CLOCK_50, waveTableSample1);
//WaveTable2Rom waveTable2Rom(waveTableIndex, CLOCK_50, waveTableSample2);

//SampleMixer sampleMixer(waveTableSample0, waveTableSample1, waveTableSample2, modulation, renderedSample);

always @(posedge CLOCK_50)
begin
	i2sCount <= i2sCount + 1'b1;
	
	if (i2sCount == i2sTicks)
		begin
			i2sCount <= 1'b0;
			
			i2sBitClock <= ~i2sBitClock;
			
			if (i2sBitClock == 1'b1)
				begin
					if (isSoundPlaying)
						i2sSoundData <= renderedSample[bitCount +: 1];
					else
						i2sSoundData <= 1'b0;
	
					if (bitCount == 0)
						begin
							i2sLeftRightSelect <= ~i2sLeftRightSelect;
							bitCount <= 15;
							
							if (i2sLeftRightSelect == 1'b1)
								begin
									waveTableIndex <= sampleIndex;
									modulation <= modulationValue;
									isSoundPlaying <= isSamplePlaying;
								end
						end
					else
						bitCount <= bitCount - 1'b1;
				end
		end
		
	noteSampleCount <= noteSampleCount + 1'b1;
	
	if (noteSampleCount >= noteSampleTicks)
		begin
			noteSampleCount <= 1'b0;
			sampleIndex <= isSamplePlaying ? sampleIndex + 1'b1 : 1'b0;
					
			if (isNoteOn == 1'b1)
				isSamplePlaying <= 1'b1;	
			else if (sampleIndex == 1'b0)
				isSamplePlaying <= 1'b0;
		end
end

endmodule

// ============================================================================
// Copyright (c) 2012 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altrea Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL or Verilog source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//
//
//
//                     web: http://www.terasic.com/
//                     email: support@terasic.com
//
// ============================================================================
//
// Major Functions:KEY triggle
//
// ============================================================================
//
// Revision History :
// ============================================================================
//   Ver  :| Author             :| Mod. Date :| Changes Made:
//   V1.0 :| Allen Wang         :| 03/25/10  :| Initial Revision
// ============================================================================



//`define  OUT_BIT  9

module keytr(
	key0,
	rst_n,
	clock,
	
	ON,				
	KEY0_EDGE,
	counter	
	);

//=======================================================
//  PORT declarations
//=======================================================			 
input			key0;
input			rst_n;
input			clock;

output			ON;
output			KEY0_EDGE;
output	[9:0]	counter;

reg     [9:0]  counter;
//reg              KEYON;
//wire ON=((counter[`OUT_BIT]==1) && (key==0))?0:1; 
/*/=============================================================================
// Structural coding
//=============================================================================
always @(negedge ON or posedge clock) 
	begin
		if (!ON)
			begin
				counter=0;
			end 
		else if (counter[`OUT_BIT]==0)
				begin
					counter=counter+1;
				end	
	end

always @(posedge clock) 
	begin
		if  ((counter>=1) && (counter <5))
			begin
				KEYON=0;
			end
		else begin	
				KEYON=1;
			 end
	end*/

///debounce starts

reg		[3:0]	flag_temp;
reg				flag;
reg		[15:0]	delay;
reg				D1;
reg 			D2;
wire			falling_edge;


//falling edge detect,
always@(negedge clock)
begin
  if (flag)
  begin 
     flag_temp<={key0, flag_temp[3:1]};
  end 
end
assign falling_edge = (flag_temp==4'b0011) ? 1'b1 : 1'b0;


////////////
always@(posedge clock,negedge rst_n)
begin
  if (!rst_n)
     flag <= 1'b1;
  else if (delay == 15'd4096)////modify the value here for a better debounce effect when using a high clock frequency;
     flag <= 1'b1;
  else if (falling_edge)
     flag <= 1'b0;
end



//
always@(posedge clock)
begin
  if (!key0)
     delay <= delay+1;
  else
     delay <= 15'd0;
end



///debounce over!
/////////////////////////////////////////
///////////?????
always@(negedge clock)
begin
  D1 <= flag;
  D2 <= D1;
end
assign KEY0_EDGE = (D1 | !D2);

endmodule	
	
// ============================================================================
// Copyright (c) 2012 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altrea Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL or Verilog source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//
//
//
//                     web: http://www.terasic.com/
//                     email: support@terasic.com
//
// ============================================================================
//
// Major Functions:i2c controller
//
// ============================================================================
//
// Revision History :
// ============================================================================
//   Ver  :| Author              :| Mod. Date :| Changes Made:
//   V1.0 :| Allen Wang          :| 03/25/10  :|      Initial Revision
//   V3.0 :| Young               :| 01/05/10  :|  vision 12.1
// ============================================================================
module i2c (
			 CLOCK,
			 I2C_SCLK,		//I2C CLOCK
			 I2C_SDAT,		//I2C DATA
			 I2C_DATA,		//DATA:[SLAVE_ADDR,SUB_ADDR,DATA]
			 GO,      		//GO transfor
			 END,    	    //END transfor 
			 W_R,     		//W_R
			 ACK,     	    //ACK
			 RESET,
			 //TEST
			 SD_COUNTER,
			 SDO
		   	);

//=======================================================
//  PORT declarations
//=======================================================
			
	input 			 CLOCK;
	input 			 [23:0]I2C_DATA;	
	input 			 GO;
	input  			 RESET;	
	input  			 W_R;
	
 	inout  			 I2C_SDAT;
 		
	output 			 I2C_SCLK;
	output			 END;	
	output 			 ACK;

//TEST
	output	[5:0]	 SD_COUNTER;
	output 			 SDO;


	reg 			 SDO;
	reg 			 SCLK;
	reg 			 END;
	reg 	[23:0]	 SD;
	reg 	[5:0]	 SD_COUNTER;

wire I2C_SCLK = SCLK | ( ((SD_COUNTER >= 4) & (SD_COUNTER <= 30))? ~CLOCK :0 );
wire I2C_SDAT = SDO?1'bz:0 ;

reg ACK1,ACK2,ACK3;
wire ACK = ACK1 | ACK2 | ACK3;

//=============================================================================
// Structural coding
//=============================================================================

//==============================I2C COUNTER====================================
always @(negedge RESET or posedge CLOCK ) 
	begin
		if (!RESET)
			begin
				SD_COUNTER = 6'b111111;
			end
		else begin
				if (GO == 0)
					begin
						SD_COUNTER = 0;
					end
				else begin
						if (SD_COUNTER < 6'b111111)
							begin
								SD_COUNTER = SD_COUNTER+1;
							end	
					 end		
			 end
	end
//==============================I2C COUNTER====================================

always @(negedge RESET or  posedge CLOCK ) 
	begin
		if (!RESET) 
			begin 
				SCLK = 1;
				SDO  = 1; 
				ACK1 = 0;
				ACK2 = 0;
				ACK3 = 0; 
				END  = 1; 
			end
		else
			case (SD_COUNTER)
					6'd0  : begin 
								ACK1 = 0 ;
								ACK2 = 0 ;
								ACK3 = 0 ; 
								END  = 0 ; 
								SDO  =1  ; 
								SCLK =1  ;
							end
					//=========start===========
					6'd1  : begin 
								SD  = I2C_DATA;
								SDO = 0;
							end
							
					6'd2  : 	SCLK = 0;
					//======SLAVE ADDR=========
					6'd3  : 	SDO = SD[23];
					6'd4  : 	SDO = SD[22];
					6'd5  : 	SDO = SD[21];
					6'd6  : 	SDO = SD[20];
					6'd7  : 	SDO = SD[19];
					6'd8  : 	SDO = SD[18];
					6'd9  :	    SDO	= SD[17];
					6'd10 : 	SDO = SD[16];	
					6'd11 : 	SDO = 1'b1;//ACK

					//========SUB ADDR==========
					6'd12  : begin 
								SDO  = SD[15]; 
								ACK1 = I2C_SDAT; 
							 end
					6'd13  : 	SDO = SD[14];
					6'd14  : 	SDO = SD[13];
					6'd15  : 	SDO = SD[12];
					6'd16  : 	SDO = SD[11];
					6'd17  : 	SDO = SD[10];
					6'd18  : 	SDO = SD[9];
					6'd19  : 	SDO = SD[8];	
					6'd20  : 	SDO = 1'b1;//ACK

					//===========DATA============
					6'd21  : begin 
								SDO  = SD[7]; 
								ACK2 = I2C_SDAT; 
							 end
					6'd22  : 	SDO = SD[6];
					6'd23  : 	SDO = SD[5];
					6'd24  : 	SDO = SD[4];
					6'd25  : 	SDO = SD[3];
					6'd26  : 	SDO = SD[2];
					6'd27  : 	SDO = SD[1];
					6'd28  : 	SDO = SD[0];	
					6'd29  : 	SDO = 1'b1;//ACK

	
					//stop
					6'd30 : begin 
								SDO  = 1'b0;	
								SCLK = 1'b0; 
								ACK3 = I2C_SDAT; 
							end	
					6'd31 : 	SCLK = 1'b1; 
					6'd32 : begin 
								SDO = 1'b1; 
								END = 1; 
							end 

			endcase
	end
	
endmodule

// ============================================================================
// Copyright (c) 2012 by Terasic Technologies Inc.
// ============================================================================
//
// Permission:
//
//   Terasic grants permission to use and modify this code for use
//   in synthesis for all Terasic Development Boards and Altrea Development 
//   Kits made by Terasic.  Other use of this code, including the selling 
//   ,duplication, or modification of any portion is strictly prohibited.
//
// Disclaimer:
//
//   This VHDL or Verilog source code is intended as a design reference
//   which illustrates how these types of functions can be implemented.
//   It is the user's responsibility to verify their design for
//   consistency and functionality through the use of formal
//   verification methods.  Terasic provides no warranty regarding the use 
//   or functionality of this code.
//
// ============================================================================
//           
//  Terasic Technologies Inc
//  9F., No.176, Sec.2, Gongdao 5th Rd, East Dist, Hsinchu City, 30070. Taiwan
//
//
//
//                     web: http://www.terasic.com/
//                     email: support@terasic.com
//
// ============================================================================
//
// Major Functions: I2C output data
//
// ============================================================================
//
// Revision History :
// ============================================================================
//   Ver  :| Author             :| Mod. Date :| Changes Made:
//   V1.0 :| Allen Wang         :| 03/24/10  :| Initial Revision
//   V3.0 :| Young       		  :| 01/05/13  :| version 12.1
// ============================================================================
`define rom_size 6'd8

module CLOCK_500(
	CLOCK,
	rst_n,
	END,
	KEY0_EDGE,
	
	DATA,
	GO,
	level_vol,				  
	CLOCK_500,				  
	CLOCK_2
	);
//=======================================================
//  PORT declarations
//=======================================================                
input  		 	CLOCK;
input 		 	rst_n;
input 		 	END;
input 		 	KEY0_EDGE;

output 	[23:0]	DATA;
output 			GO;
output	[3:0] 	level_vol;
output		    CLOCK_500;
output 			CLOCK_2;


reg  	[10:0]	COUNTER_500;
reg  	[15:0]	ROM[`rom_size:0];
reg  	[15:0]	DATA_A;
reg  	[5:0]	address;




wire  CLOCK_500 = COUNTER_500[9];
wire  CLOCK_2 	= COUNTER_500[1];

wire [23:0]DATA = {8'h34, DATA_A};		//slave address + sub_address + register_data
wire  GO = ((address <= `rom_size) && (END == 1)) ? COUNTER_500[10] : 1;
//=============================================================================
// Structural coding
//=============================================================================

always @(posedge CLOCK ) 
begin
	COUNTER_500=COUNTER_500+1;
end


always @(negedge KEY0_EDGE or posedge END) 
begin
	if (!KEY0_EDGE)
	begin
		address=0;
	end
	else if (address <= `rom_size)
	begin
		address=address+1;
	end
end

reg		[4:0]	vol;
wire	[6:0]	volume;

always @(negedge KEY0_EDGE or negedge rst_n) 
begin
	if(!rst_n)
		vol = 5'd31;
	else if(vol == 5'd4)
		vol = 5'd31;
	else if(!KEY0_EDGE)
		vol = vol - 3;
end

//the volume level, level 0 to level 9,
//the higher the level, the greater the sound
assign level_vol = (vol - 4) / 3;
assign volume = vol + 96;


always @(posedge END) 
begin
	ROM[0] = 16'h0c00;	    			 	//power down
	ROM[1] = 16'h0ec2;	   		    	 	//master
	ROM[2] = 16'h0838;	    			 	//sound select
	
	ROM[3] = 16'h1000;						//mclk
	
	ROM[4] = 16'h0017;						//
	ROM[5] = 16'h0217;					 	//
	ROM[6] = {8'h04,1'b0,volume[6:0]};		//left channel headphone output volume
	ROM[7] = {8'h06,1'b0,volume[6:0]};		//right channel headphone output volume
	
	//ROM[4]= 16'h1e00;		             	//reset	
	ROM[`rom_size] = 16'h1201;           	//active
	DATA_A = ROM[address];
end


endmodule

module  HEX(
input	[3:0]	hex,
output	[6:0]	hex_fps
);


assign hex_fps	=	(hex == 4'd0) ? 7'h40: //0
					(hex == 4'd1) ? 7'h79: //1
					(hex == 4'd2) ? 7'h24: //2
					(hex == 4'd3) ? 7'h30: //3
					(hex == 4'd4) ? 7'h19: //4        
					(hex == 4'd5) ? 7'h12: //5
					(hex == 4'd6) ? 7'h02: //6
					(hex == 4'd7) ? 7'h78: //7
					(hex == 4'd8) ? 7'h00: //8
									7'h10; //9

endmodule 